module counter(input clk,
              input rstn,
              input clear,
              input incr,
              output reg [2:0] count);
  
  
  
  
  
  always @(posedge clk,negedge rstn)
    begin
      if(!rstn)
        count<='b0;
      else if(clear)
        count<='b0;
      else
        count<=count+incr;
    end
  
  
endmodule
