module tb_shift_reg;
  reg clk;
  reg rstn;
  reg shift_en;
  reg data_in;
  wire [4:0] data_out;
  
  shift_reg_n #(.n(5)) dut1(.clk(clk),
                           .rstn(rstn),
                           .data_in(data_in),
                           .shift_en(shift_en),
                           .data_out(data_out));
  
  
  initial begin
    
    $dumpfile("dump.vcd");
    $dumpvars(1);
    
    clk=1;
    rstn=0;
    shift_en=0;
    data_in='b0;
    
    repeat (5) begin
      
    #10 rstn=1;
      
    shift_en=1;
    data_in=1;
      
    #10 data_in=1;
    #10 data_in=1;
    #10 data_in=1;
    #10 data_in=1;
    #10 rstn=0;
    shift_en=0;
      
    end

    
  end
  
  always #5 clk=~clk;
                
  initial #300 $finish;
  
  
endmodule
